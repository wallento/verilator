module t;

endmodule