module timescalemod;

endmodule